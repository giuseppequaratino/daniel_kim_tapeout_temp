// OpenRAM SRAM model
// Words: 4096 (2^12)
// Word size: 32
// Write size: 8

module sram(
`ifdef USE_POWER_PINS
    vccd1,
    vssd1,
`endif
// Port 0: RW
    clk0,csb0,web0,wmask0,addr0,din0,dout0, //wmask not used
// Port 1: R
    clk1,csb1,addr1,dout1,
// Port 2: R
    clk2,csb2,addr2,dout2
  );
	//1280x720 --> 80x45 blocks = 3600 blocks -->4096 = 2^12
  parameter NUM_WMASKS = 4 ;
  parameter DATA_WIDTH = 2048 ;//16x16x8 = 2048
  parameter ADDR_WIDTH = 12 ;
  parameter RAM_DEPTH = 1 << ADDR_WIDTH;
  // FIXME: This delay is arbitrary.
  parameter DELAY = 3 ;
  parameter VERBOSE = 1 ; //Set to 0 to only display warnings
  parameter T_HOLD = 1 ; //Delay to hold dout value after posedge. Value is arbitrary

`ifdef USE_POWER_PINS
    inout vccd1;
    inout vssd1;
`endif
  input  clk0; // clock
  input   csb0; // active low chip select
  input  web0; // active low write control
  input [NUM_WMASKS-1:0]   wmask0; // write mask
  input [ADDR_WIDTH-1:0]  addr0;
  input [DATA_WIDTH-1:0]  din0;
  output [DATA_WIDTH-1:0] dout0;
  input  clk1; // clock
  input   csb1; // active low chip select
  input [ADDR_WIDTH-1:0]  addr1;
  output [DATA_WIDTH-1:0] dout1;

  input clk2;
  input csb2;
  input [ADDR_WIDTH-1:0] addr2;
  output [DATA_WIDTH-1:0] dout2;





  reg  csb0_reg;
  reg  web0_reg;
  reg [NUM_WMASKS-1:0]   wmask0_reg;
  reg [ADDR_WIDTH-1:0]  addr0_reg;
  reg [DATA_WIDTH-1:0]  din0_reg;
  reg [DATA_WIDTH-1:0]  dout0;

  // All inputs are registers
  always @(posedge clk0)
  begin
    csb0_reg = csb0;
    web0_reg = web0;
    wmask0_reg = wmask0;
    addr0_reg = addr0;
    din0_reg = din0;
    #(T_HOLD) dout0 = 2048'bx;
    if ( !csb0_reg && web0_reg && VERBOSE ) 
      $display($time," Reading %m addr0=%d dout0=%b",addr0_reg,mem[addr0_reg]);
    if ( !csb0_reg && !web0_reg && VERBOSE )
      $display($time," Writing %m addr0=%d din0=%h wmask0=%b",addr0_reg,din0_reg,wmask0_reg);
  end

  reg  csb1_reg;
  reg [ADDR_WIDTH-1:0]  addr1_reg;
  reg [DATA_WIDTH-1:0]  dout1;


  reg  csb2_reg;
  reg [ADDR_WIDTH-1:0]  addr2_reg;
  reg [DATA_WIDTH-1:0]  dout2;

  // All inputs are registers
  always @(posedge clk1)
  begin
    csb1_reg = csb1;
    addr1_reg = addr1;
    if (!csb0 && !web0 && !csb1 && (addr0 == addr1))
         $display($time," WARNING: Writing and reading addr0=%d and addr1=%d simultaneously!",addr0,addr1);
    #(T_HOLD) dout1 = 2048'bx;
    if ( !csb1_reg && VERBOSE ) 
      $display($time," Reading %m addr1=%d dout1=%b",addr1_reg,mem[addr1_reg]);
  end

  always @(posedge clk2) begin
    csb2_reg = csb2;
    addr2_reg = addr2;
    if ( !csb2_reg && VERBOSE ) 
      $display($time," Reading %m addr1=%d dout1=%b",addr2_reg,mem[addr2_reg]);
  end


reg [DATA_WIDTH-1:0]    mem [0:RAM_DEPTH-1];

  // Memory Write Block Port 0
  // Write Operation : When web0 = 0, csb0 = 0
  always @ (negedge clk0)
  begin : MEM_WRITE0
    if ( !csb0_reg && !web0_reg ) begin
            mem[addr0_reg] = din0_reg;
    end
  end

  // Memory Read Block Port 0
  // Read Operation : When web0 = 1, csb0 = 0
  always @ (negedge clk0)
  begin : MEM_READ0
    if (!csb0_reg && web0_reg)
       dout0 <= #(DELAY) mem[addr0_reg];
  end

  // Memory Read Block Port 1
  // Read Operation : When web1 = 1, csb1 = 0
  always @ (negedge clk1)
  begin : MEM_READ1
    if (!csb1_reg)
       dout1 <= #(DELAY) mem[addr1_reg];
  end

  // Memory Read Block Port 1
  // Read Operation : When web1 = 1, csb1 = 0
  always @ (negedge clk2)
  begin : MEM_READ2
    if (!csb2_reg)
       dout2 <= #(DELAY) mem[addr2_reg];
  end

endmodule
